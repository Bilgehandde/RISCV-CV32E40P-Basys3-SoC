`timescale 1ns / 1ps

module simple_ram #(
    parameter SIZE_WORDS = 1024 // 1024 kelime = 4KB Haf�za
)(
    input  logic        clk,
    input  logic        rst_n,
    
    // ��lemciden gelen sinyaller
    input  logic        req_i,       // "Veri istiyorum" sinyali
    input  logic        we_i,        // "Yazma yap�cam" sinyali (0 ise Okuma)
    input  logic [31:0] addr_i,      // "Hangi adresteki veri?"
    input  logic [31:0] wdata_i,     // Yaz�lacak veri
    input  logic [3:0]  be_i,        // Byte Enable (Hangi byte'lar� yazal�m?)
    
    // ��lemciye giden sinyaller
    output logic [31:0] rdata_o,     // Okunan veri
    output logic        rvalid_o     // "Veri haz�r" sinyali
);

    // 1. Haf�za Dizisi (As�l Depo)
    // 32 bit geni�li�inde, 1024 sat�rl�k bir tablo
    logic [31:0] mem [0:SIZE_WORDS-1];

    // 2. Ba�lang��ta ��ini Doldur (Yaz�l�m� Y�kle)
    initial begin
        // program.hex dosyas�n� okuyup haf�zaya yazar
        // Bu dosyan�n projenin sim�lasyon klas�r�nde olmas� laz�m!
        $readmemh("program.hex", mem);
    end

    // 3. Okuma ve Yazma Mant���
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rdata_o  <= 32'h0;
            rvalid_o <= 1'b0;
        end else begin
            // Varsay�lan olarak valid 0 olsun
            rvalid_o <= 1'b0;

            if (req_i) begin
                // E�er istek varsa 1 �evrim sonra cevap ver (Synchronous RAM)
                rvalid_o <= 1'b1;

                if (we_i) begin
                    // --- YAZMA ��LEM� ---
                    // RISC-V adresleri byte bazl�d�r (0, 4, 8...). 
                    // Ama bizim dizimiz word bazl� (0, 1, 2...). 
                    // O y�zden adresi 4'e b�l�yoruz (addr_i >> 2).
                    if (be_i[0]) mem[addr_i[31:2]][7:0]   <= wdata_i[7:0];
                    if (be_i[1]) mem[addr_i[31:2]][15:8]  <= wdata_i[15:8];
                    if (be_i[2]) mem[addr_i[31:2]][23:16] <= wdata_i[23:16];
                    if (be_i[3]) mem[addr_i[31:2]][31:24] <= wdata_i[31:24];
                end else begin
                    // --- OKUMA ��LEM� ---
                    rdata_o <= mem[addr_i[31:2]];
                end
            end
        end
    end

endmodule